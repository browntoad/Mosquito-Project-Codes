`timescale	1ns/1ns
module top_tb;

    //	Internal Regs and Nets
    reg	 clk;
    reg	 rst;
    reg [15:0] din;
    wire in_en;
    wire is_mosq;

    localparam N = 5000;
    // localparam N = 24000;    
    integer tp;

    reg signed [15:0] in_mem[0:N-1];

    assign in_en = ~rst;

    top DUT (
        .din(din),
        .in_en(in_en),
        .clk(clk),
        .rst(rst),
        .is_mosq(is_mosq)
    );

//----------------------------------------------------------------------
//	Clock and Reset
//----------------------------------------------------------------------
    initial begin
        clk <= 1;
        rst <= 1;
        forever #5 clk <= ~clk;
    end

    // initial begin
    //     $fsdbDumpfile("top.fsdb");
    //     $fsdbDumpvars("+mda");
    // end

//----------------------------------------------------------------------
//	Tasks
//----------------------------------------------------------------------

    task GenerateInputWave;
        input[80*8:1] filename;
        input[63:0] case_idx;
        integer n;
    begin
        $readmemh(filename, in_mem);

        @(posedge clk);
        rst <= 0;

        for (n = 0; n < N; n = n + 1) begin
            din <= (in_mem[n]/16);
            @(posedge clk);
        end
        
        din <= 0;

        repeat(500) @(posedge clk);
        $display("Test case %d: is_mosq = %d", case_idx, is_mosq);
        rst <= 1;
        tp = tp + is_mosq;
        repeat(10) @(posedge clk);
    end
    endtask

    initial begin
        repeat(10) @(posedge clk);
        tp = 0;
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_001.txt", 000);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_002.txt", 001);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_003.txt", 002);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_004.txt", 003);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_005.txt", 004);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_006.txt", 005);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_007.txt", 006);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_008.txt", 007);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_009.txt", 008);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_010.txt", 009);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_011.txt", 010);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_012.txt", 011);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_013.txt", 012);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_014.txt", 013);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_015.txt", 014);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_016.txt", 015);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_017.txt", 016);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_018.txt", 017);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_019.txt", 018);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_020.txt", 019);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_021.txt", 020);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_022.txt", 021);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_023.txt", 022);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_024.txt", 023);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_025.txt", 024);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_026.txt", 025);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_027.txt", 026);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_028.txt", 027);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_029.txt", 028);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_030.txt", 029);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_031.txt", 030);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_032.txt", 031);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_033.txt", 032);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_034.txt", 033);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_035.txt", 034);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_036.txt", 035);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_037.txt", 036);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_038.txt", 037);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_039.txt", 038);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_040.txt", 039);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_041.txt", 040);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_042.txt", 041);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_043.txt", 042);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_044.txt", 043);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_045.txt", 044);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_046.txt", 045);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_047.txt", 046);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_048.txt", 047);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_049.txt", 048);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_050.txt", 049);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_051.txt", 050);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_052.txt", 051);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_053.txt", 052);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_054.txt", 053);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_055.txt", 054);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_056.txt", 055);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_057.txt", 056);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_058.txt", 057);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_059.txt", 058);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_060.txt", 059);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_061.txt", 060);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_062.txt", 061);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_063.txt", 062);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_064.txt", 063);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_065.txt", 064);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_066.txt", 065);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_067.txt", 066);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_068.txt", 067);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_069.txt", 068);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_070.txt", 069);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_071.txt", 070);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_072.txt", 071);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_073.txt", 072);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_074.txt", 073);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_075.txt", 074);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_076.txt", 075);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_077.txt", 076);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_078.txt", 077);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_079.txt", 078);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_080.txt", 079);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_081.txt", 080);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_082.txt", 081);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_083.txt", 082);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_084.txt", 083);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_085.txt", 084);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_086.txt", 085);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_087.txt", 086);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_088.txt", 087);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_089.txt", 088);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_090.txt", 089);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_091.txt", 090);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_092.txt", 091);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_093.txt", 092);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_094.txt", 093);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_095.txt", 094);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_096.txt", 095);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_097.txt", 096);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_098.txt", 097);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_099.txt", 098);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_100.txt", 099); 
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_101.txt", 100);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_102.txt", 101);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_103.txt", 102);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_104.txt", 103);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_105.txt", 104);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_106.txt", 105);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_107.txt", 106);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_108.txt", 107);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_109.txt", 108);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_110.txt", 109);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_111.txt", 110);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_112.txt", 111);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_113.txt", 112);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_114.txt", 113);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_115.txt", 114);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_116.txt", 115);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_117.txt", 116);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_118.txt", 117);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_119.txt", 118);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_120.txt", 119);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_121.txt", 120);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_122.txt", 121);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_123.txt", 122);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_124.txt", 123);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_125.txt", 124);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_126.txt", 125);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_127.txt", 126);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_128.txt", 127);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_129.txt", 128);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_130.txt", 129);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_131.txt", 130);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_132.txt", 131);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_133.txt", 132);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_134.txt", 133);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_135.txt", 134);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_136.txt", 135);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_137.txt", 136);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_138.txt", 137);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_139.txt", 138);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_140.txt", 139);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_141.txt", 140);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_142.txt", 141);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_143.txt", 142);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_144.txt", 143);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_145.txt", 144);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_146.txt", 145);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_147.txt", 146);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_148.txt", 147);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_149.txt", 148);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_150.txt", 149); 
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_151.txt", 150);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_152.txt", 151);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_153.txt", 152);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_154.txt", 153);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_155.txt", 154);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_156.txt", 155);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_157.txt", 156);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_158.txt", 157);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_159.txt", 158);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_160.txt", 159);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_161.txt", 160);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_162.txt", 161);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_163.txt", 162);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_164.txt", 163);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_165.txt", 164);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_166.txt", 165);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_167.txt", 166);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_168.txt", 167);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_169.txt", 168);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_170.txt", 169);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_171.txt", 170);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_172.txt", 171);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_173.txt", 172);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_174.txt", 173);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_175.txt", 174);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_176.txt", 175);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_177.txt", 176);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_178.txt", 177);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_179.txt", 178);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_180.txt", 179);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_181.txt", 180);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_182.txt", 181);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_183.txt", 182);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_184.txt", 183);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_185.txt", 184);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_186.txt", 185);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_187.txt", 186);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_188.txt", 187);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_189.txt", 188);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_190.txt", 189);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_191.txt", 190);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_192.txt", 191);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_193.txt", 192);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_194.txt", 193);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_195.txt", 194);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_196.txt", 195);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_197.txt", 196);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_198.txt", 197);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_199.txt", 198);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_200.txt", 199); 
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_201.txt", 200);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_202.txt", 201);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_203.txt", 202);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_204.txt", 203);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_205.txt", 204);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_206.txt", 205);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_207.txt", 206);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_208.txt", 207);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_209.txt", 208);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_210.txt", 209);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_211.txt", 210);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_212.txt", 211);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_213.txt", 212);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_214.txt", 213);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_215.txt", 214);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_216.txt", 215);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_217.txt", 216);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_218.txt", 217);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_219.txt", 218);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_220.txt", 219);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_221.txt", 220);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_222.txt", 221);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_223.txt", 222);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_224.txt", 223);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_225.txt", 224);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_226.txt", 225);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_227.txt", 226);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_228.txt", 227);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_229.txt", 228);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_230.txt", 229);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_231.txt", 230);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_232.txt", 231);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_233.txt", 232);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_234.txt", 233);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_235.txt", 234);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_236.txt", 235);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_237.txt", 236);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_238.txt", 237);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_239.txt", 238);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_240.txt", 239);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_241.txt", 240);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_242.txt", 241);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_243.txt", 242);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_244.txt", 243);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_245.txt", 244);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_246.txt", 245);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_247.txt", 246);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_248.txt", 247);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_249.txt", 248);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_250.txt", 249); 
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_251.txt", 250);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_252.txt", 251);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_253.txt", 252);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_254.txt", 253);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_255.txt", 254);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_256.txt", 255);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_257.txt", 256);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_258.txt", 257);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_259.txt", 258);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_260.txt", 259);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_261.txt", 260);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_262.txt", 261);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_263.txt", 262);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_264.txt", 263);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_265.txt", 264);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_266.txt", 265);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_267.txt", 266);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_268.txt", 267);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_269.txt", 268);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_270.txt", 269);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_271.txt", 270);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_272.txt", 271);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_273.txt", 272);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_274.txt", 273);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_275.txt", 274);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_276.txt", 275);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_277.txt", 276);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_278.txt", 277);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_279.txt", 278);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_280.txt", 279);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_281.txt", 280);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_282.txt", 281);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_283.txt", 282);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_284.txt", 283);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_285.txt", 284);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_286.txt", 285);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_287.txt", 286);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_288.txt", 287);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_289.txt", 288);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_290.txt", 289);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_291.txt", 290);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_292.txt", 291);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_293.txt", 292);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_294.txt", 293);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_295.txt", 294);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_296.txt", 295);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_297.txt", 296);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_298.txt", 297);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_299.txt", 298);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_300.txt", 299); 
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_301.txt", 300);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_302.txt", 301);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_303.txt", 302);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_304.txt", 303);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_305.txt", 304);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_306.txt", 305);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_307.txt", 306);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_308.txt", 307);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_309.txt", 308);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_310.txt", 309);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_311.txt", 310);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_312.txt", 311);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_313.txt", 312);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_314.txt", 313);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_315.txt", 314);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_316.txt", 315);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_317.txt", 316);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_318.txt", 317);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_319.txt", 318);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_320.txt", 319);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_321.txt", 320);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_322.txt", 321);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_323.txt", 322);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_324.txt", 323);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_325.txt", 324);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_326.txt", 325);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_327.txt", 326);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_328.txt", 327);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_329.txt", 328);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_330.txt", 329);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_331.txt", 330);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_332.txt", 331);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_333.txt", 332);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_334.txt", 333);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_335.txt", 334);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_336.txt", 335);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_337.txt", 336);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_338.txt", 337);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_339.txt", 338);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_340.txt", 339);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_341.txt", 340);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_342.txt", 341);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_343.txt", 342);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_344.txt", 343);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_345.txt", 344);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_346.txt", 345);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_347.txt", 346);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_348.txt", 347);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_349.txt", 348);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_350.txt", 349); 
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_351.txt", 350);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_352.txt", 351);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_353.txt", 352);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_354.txt", 353);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_355.txt", 354);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_356.txt", 355);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_357.txt", 356);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_358.txt", 357);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_359.txt", 358);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_360.txt", 359);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_361.txt", 360);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_362.txt", 361);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_363.txt", 362);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_364.txt", 363);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_365.txt", 364);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_366.txt", 365);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_367.txt", 366);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_368.txt", 367);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_369.txt", 368);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_370.txt", 369);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_371.txt", 370);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_372.txt", 371);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_373.txt", 372);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_374.txt", 373);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_375.txt", 374);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_376.txt", 375);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_377.txt", 376);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_378.txt", 377);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_379.txt", 378);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_380.txt", 379);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_381.txt", 380);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_382.txt", 381);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_383.txt", 382);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_384.txt", 383);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_385.txt", 384);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_386.txt", 385);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_387.txt", 386);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_388.txt", 387);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_389.txt", 388);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_390.txt", 389);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_391.txt", 390);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_392.txt", 391);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_393.txt", 392);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_394.txt", 393);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_395.txt", 394);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_396.txt", 395);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_397.txt", 396);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_398.txt", 397);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_399.txt", 398);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_400.txt", 399); 
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_401.txt", 400);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_402.txt", 401);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_403.txt", 402);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_404.txt", 403);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_405.txt", 404);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_406.txt", 405);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_407.txt", 406);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_408.txt", 407);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_409.txt", 408);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_410.txt", 409);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_411.txt", 410);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_412.txt", 411);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_413.txt", 412);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_414.txt", 413);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_415.txt", 414);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_416.txt", 415);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_417.txt", 416);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_418.txt", 417);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_419.txt", 418);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_420.txt", 419);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_421.txt", 420);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_422.txt", 421);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_423.txt", 422);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_424.txt", 423);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_425.txt", 424);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_426.txt", 425);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_427.txt", 426);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_428.txt", 427);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_429.txt", 428);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_430.txt", 429);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_431.txt", 430);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_432.txt", 431);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_433.txt", 432);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_434.txt", 433);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_435.txt", 434);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_436.txt", 435);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_437.txt", 436);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_438.txt", 437);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_439.txt", 438);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_440.txt", 439);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_441.txt", 440);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_442.txt", 441);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_443.txt", 442);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_444.txt", 443);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_445.txt", 444);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_446.txt", 445);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_447.txt", 446);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_448.txt", 447);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_449.txt", 448);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_450.txt", 449); 
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_451.txt", 450);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_452.txt", 451);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_453.txt", 452);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_454.txt", 453);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_455.txt", 454);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_456.txt", 455);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_457.txt", 456);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_458.txt", 457);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_459.txt", 458);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_460.txt", 459);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_461.txt", 460);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_462.txt", 461);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_463.txt", 462);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_464.txt", 463);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_465.txt", 464);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_466.txt", 465);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_467.txt", 466);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_468.txt", 467);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_469.txt", 468);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_470.txt", 469);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_471.txt", 470);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_472.txt", 471);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_473.txt", 472);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_474.txt", 473);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_475.txt", 474);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_476.txt", 475);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_477.txt", 476);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_478.txt", 477);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_479.txt", 478);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_480.txt", 479);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_481.txt", 480);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_482.txt", 481);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_483.txt", 482);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_484.txt", 483);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_485.txt", 484);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_486.txt", 485);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_487.txt", 486);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_488.txt", 487);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_489.txt", 488);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_490.txt", 489);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_491.txt", 490);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_492.txt", 491);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_493.txt", 492);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_494.txt", 493);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_495.txt", 494);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_496.txt", 495);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_497.txt", 496);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_498.txt", 497);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_499.txt", 498);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_500.txt", 499); 
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_501.txt", 500);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_502.txt", 501);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_503.txt", 502);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_504.txt", 503);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_505.txt", 504);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_506.txt", 505);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_507.txt", 506);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_508.txt", 507);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_509.txt", 508);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_510.txt", 509);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_511.txt", 510);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_512.txt", 511);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_513.txt", 512);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_514.txt", 513);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_515.txt", 514);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_516.txt", 515);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_517.txt", 516);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_518.txt", 517);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_519.txt", 518);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_520.txt", 519);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_521.txt", 520);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_522.txt", 521);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_523.txt", 522);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_524.txt", 523);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_525.txt", 524);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_526.txt", 525);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_527.txt", 526);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_528.txt", 527);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_529.txt", 528);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_530.txt", 529);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_531.txt", 530);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_532.txt", 531);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_533.txt", 532);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_534.txt", 533);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_535.txt", 534);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_536.txt", 535);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_537.txt", 536);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_538.txt", 537);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_539.txt", 538);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_540.txt", 539);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_541.txt", 540);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_542.txt", 541);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_543.txt", 542);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_544.txt", 543);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_545.txt", 544);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_546.txt", 545);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_547.txt", 546);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_548.txt", 547);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_549.txt", 548);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_550.txt", 549); 
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_551.txt", 550);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_552.txt", 551);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_553.txt", 552);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_554.txt", 553);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_555.txt", 554);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_556.txt", 555);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_557.txt", 556);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_558.txt", 557);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_559.txt", 558);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_560.txt", 559);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_561.txt", 560);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_562.txt", 561);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_563.txt", 562);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_564.txt", 563);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_565.txt", 564);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_566.txt", 565);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_567.txt", 566);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_568.txt", 567);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_569.txt", 568);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_570.txt", 569);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_571.txt", 570);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_572.txt", 571);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_573.txt", 572);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_574.txt", 573);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_575.txt", 574);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_576.txt", 575);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_577.txt", 576);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_578.txt", 577);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_579.txt", 578);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_580.txt", 579);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_581.txt", 580);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_582.txt", 581);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_583.txt", 582);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_584.txt", 583);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_585.txt", 584);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_586.txt", 585);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_587.txt", 586);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_588.txt", 587);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_589.txt", 588);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_590.txt", 589);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_591.txt", 590);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_592.txt", 591);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_593.txt", 592);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_594.txt", 593);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_595.txt", 594);             
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_596.txt", 595);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_597.txt", 596);    
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_598.txt", 597);
        GenerateInputWave("C:/Users/isaia/Downloads/mosq_proj/pat/mosq/mosq_599.txt", 598);
        $display("tp = %d", tp);
        $display("fp = %d", (599-tp));

        repeat(10) @(posedge clk);
        $finish;
    end

    initial begin
        repeat(20000000) @(posedge clk);
        $display("[FAILED] Simulation timed out.");
        $finish;
    end

endmodule
